`timescale 1 ps / 1 ps

module aes32_dsp_8p_func_dec (
  input  wire         CLK,  
  input  wire         RST,
  input  wire [31:00] DIN,
  input  wire [31:00] PTX,  
  input  wire [31:00] KEY,
  input  wire [03:00] TSH, // T-table shift control (shifts the output of the BRAMs)
  input  wire [07:00] BCT, // BRAM control; [7:4] choose between T0 and T2; [3:0] chooses last round's T-tables 
  input  wire         POB, // select: plaintext(HIGH) or BRAM(LOW)
  input  wire [02:00] RXR, // reset input to DSP (so data it unchanged as it passes through)
  
  output wire [31:00] DOUT
);

  // DSP48E OPMODE settings (see UG193)
  parameter C_XOR_AB = 7'b0110011;
  parameter PCIN_XOR_AB = 7'b0010011;

  reg    [31:00] bram0a_data_p, bram0b_data_p, bram1a_data_p, bram1b_data_p;
  
  wire   [31:00] dsp0a_din;
  wire   [47:00] dsp0a_pdata, dsp0b_pdata, dsp1a_pdata, dsp1b_pdata;
  wire   [31:00] bram0a_data, bram0b_data, bram1a_data, bram1b_data;
  wire   [15:00] bram0a_addr, bram0b_addr, bram1a_addr, bram1b_addr;

  assign DOUT = dsp1b_pdata[31:00];  

  // address busses for the BRAMs {0,T0/T2,LAST,DATA,00000}
  assign bram0a_addr = {1'b0, BCT[7], BCT[3], DIN[31:24], 5'd0};
  assign bram0b_addr = {1'b0, BCT[6], BCT[2], DIN[23:16], 5'd0};
  assign bram1a_addr = {1'b0, BCT[5], BCT[1], DIN[15:08], 5'd0};
  assign bram1b_addr = {1'b0, BCT[4], BCT[0], DIN[07:00], 5'd0};
  
  // for simulation
  initial begin
    bram0a_data_p = 0; bram0b_data_p = 0; bram1a_data_p = 0; bram1b_data_p = 0;
  end  

  RAMB36 #(
    .DOA_REG            (1              ), // Optional output registers on A port (0 or 1)
    .DOB_REG            (1              ), // Optional output registers on B port (0 or 1)
    .INIT_A             (36'h000000000  ), // Initial values on A output port
    .INIT_B             (36'h000000000  ), // Initial values on B output port
    .RAM_EXTENSION_A    ("NONE"         ), // "UPPER", "LOWER" or "NONE" when cascaded
    .RAM_EXTENSION_B    ("NONE"         ), // "UPPER", "LOWER" or "NONE" when cascaded
    .READ_WIDTH_A       (36             ), // Valid values are 1, 2, 4, 9, 18, or 36
    .READ_WIDTH_B       (36             ), // Valid values are 1, 2, 4, 9, 18, or 36
    .SIM_COLLISION_CHECK("NONE"         ), // Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
    .SRVAL_A            (36'h000000000  ), // Set/Reset value for A port output
    .SRVAL_B            (36'h000000000  ), // Set/Reset value for B port output
    .WRITE_MODE_A       ("READ_FIRST"   ), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
    .WRITE_MODE_B       ("READ_FIRST"   ), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
    .WRITE_WIDTH_A      (36             ), // Valid values are 1, 2, 4, 9, 18, or 36
    .WRITE_WIDTH_B      (36             ), // Valid values are 1, 2, 4, 9, 18, or 36

   // TABLE T0 (t_in)
   .INIT_00(256'h4BE30393ACFA58AB1F9D45F13BAB6BCB3A275E961A17A4C37E41655351F4A750),
   .INIT_01(256'hB562A38F26354480C52ACBD74FE5D7FCF5024C2588CC7691AD766DF62030FA55),
   .INIT_02(256'h6BD3F9C68D4697A3814CF012C32F75025DFEC0E145EA0E9825BA1B67DEB15A49),
   .INIT_03(256'h8EC9C84449E06929587421D3D4BE832D955259DABF6D7AEB15929C95038F5FE7),
   .INIT_04(256'h7DCE3AB4C920AC66F088AD17BEE14FB627B971DD99583E6BF48E797875C2896A),
   .INIT_05(256'hF9082B94FE81A01CBB6BAE84B16477E062537F4597513360E51A318263DF4A18),
   .INIT_06(256'h6655AB2AE31F8F57724B02E2AB73D323527BF8B794DE6C878F45FD1970486858),
   .INIT_07(256'hED16825C02036ABA23BFA5B2302887F2D33708A586C57B9A2FB5C203B2EB2807),
   .INIT_08(256'hC4A6FE8AD134621F0605BED565DAF4CD4E69E2A1F307F2F0A779B4928ACF1C2B),
   .INIT_09(256'hBD6E10515E719F064060EFAA0B83EC39A4F6EB75058AE132A2F355A0342E539D),
   .INIT_0A(256'h605015FF0406D46F71C45D0591548DB54DE6BD46DD3E05AE96DD063D3E218AF9),
   .INIT_0B(256'h79C8EEDBE7195B3807898B88B0E842BD67D99E77894043CCD6BDE9971998FB24),
   .INIT_0C(256'h6C5A724E1E1170AC322BED480980868300000000F8841EC97C420FE9A17C0A47),
   .INIT_0D(256'h24362E3A9B5B54D1685CA6210A0FD964362D39273DAED51E0F853856FD0EFFFB),
   .INIT_0E(256'h1C121A165A774B6961DC20A280C0C54F1B9B919EB4EE96D29357E70F0C0A67B1),
   .INIT_0F(256'h141EA9C82DB6A8B9F28BC7AD0E090D0B121B171D3C22E043C0A02AE5E293BA0A),
   .INIT_10(256'h5BFB7E3444663BC55C72F5BCF701269FA37F60FDEE99DDBBAF75074C57F11985),
   .INIT_11(256'h84C611201397224042638510D731DCCAB8E4F163B6EDFC68CB23C6DC8B432976),
   .INIT_12(256'h77C1E3D00D8652ECDCB230F31D9E2F4BC729A16DAEF93211D2BB3DF8854A247D),
   .INIT_13(256'h223390EF567D2CD8A0F03F1AA8FC8CC447E96422119448FAA970B9992BB3166C),
   .INIT_14(256'h3FADBFA4DAB78E26A57ADE28A6F581CF98D40B368CCAA2FED938D1C187494EC7),
   .INIT_15(256'h82C3AFF52E39F75E90D8B8E8F68D13C2547E46626A5FCC9B5078920D2C3A9DE4),
   .INIT_16(256'hDB3BBB7BE89C636E10187DA7C8AC993BCF2512B36FD52DA969D0937C9F5D80BE),
   .INIT_17(256'hEF15E8E621BCCF08AAFFE67EE6956E65834F9AA8EC9AB7016E5918F4CD267809),
   .INIT_18(256'h35A266C0C6A594302A3F233131A4B2AF29B07CD6EA9F09D44A6F36CEBAE79BD9),
   .INIT_19(256'h1791F62F7FCD500E41ECDAF7F104984A33A7D815E090D0B0FC82CAA6744EBC37),
   .INIT_1A(256'h4665517FC12C1FB84C6A881B9ED1B5E3E49604DFCCAA4D5443EFB04D764DD68D),
   .INIT_1B(256'h6DD64713E910563392DBD252B3671D5AFB0B412EFA877473018C355D9D5EEA04),
   .INIT_1C(256'h7A47B13CE11CE5EDB761C935CEA927EEEB133C8959F8148E37A10C7A9AD7618C),
   .INIT_1D(256'h7844DB86DF3D6F145FFDAA5B53F7CDEA73C737BF1814CE7955F2733F9CD2DF59),
   .INIT_1E(256'hFF0D9541283C498BBCE2250C161DC372C2A3405F3824342CB968C43ECAAFF381),
   .INIT_1F(256'hD0B85742486C5C74D532B6707BCB84616456C190D8B4E49C080CB3DE39A80171),
   // TABLE T0 (t_il)
   .INIT_20(256'h38000000A50000003600000030000000D50000006A0000000900000052000000),
   .INIT_21(256'hFB000000D7000000F3000000810000009E000000A300000040000000BF000000),
   .INIT_22(256'h87000000FF0000002F0000009B0000008200000039000000E30000007C000000),
   .INIT_23(256'hCB000000E9000000DE000000C400000044000000430000008E00000034000000),
   .INIT_24(256'h3D00000023000000C2000000A600000032000000940000007B00000054000000),
   .INIT_25(256'h4E000000C3000000FA000000420000000B000000950000004C000000EE000000),
   .INIT_26(256'hB200000024000000D90000002800000066000000A10000002E00000008000000),
   .INIT_27(256'h25000000D10000008B0000006D00000049000000A20000005B00000076000000),
   .INIT_28(256'h1600000098000000680000008600000064000000F6000000F800000072000000),
   .INIT_29(256'h92000000B6000000650000005D000000CC0000005C000000A4000000D4000000),
   .INIT_2A(256'hDA000000B9000000ED000000FD0000005000000048000000700000006C000000),
   .INIT_2B(256'h840000009D0000008D000000A70000005700000046000000150000005E000000),
   .INIT_2C(256'h0A000000D3000000BC0000008C00000000000000AB000000D800000090000000),
   .INIT_2D(256'h0600000045000000B3000000B80000000500000058000000E4000000F7000000),
   .INIT_2E(256'h020000000F0000003F000000CA0000008F0000001E0000002C000000D0000000),
   .INIT_2F(256'h6B0000008A000000130000000100000003000000BD000000AF000000C1000000),
   .INIT_30(256'hEA000000DC000000670000004F0000004100000011000000910000003A000000),
   .INIT_31(256'h73000000E6000000B4000000F0000000CE000000CF000000F200000097000000),
   .INIT_32(256'h8500000035000000AD000000E70000002200000074000000AC00000096000000),
   .INIT_33(256'h6E000000DF000000750000001C000000E800000037000000F9000000E2000000),
   .INIT_34(256'h89000000C5000000290000001D000000710000001A000000F100000047000000),
   .INIT_35(256'h1B000000BE00000018000000AA0000000E00000062000000B70000006F000000),
   .INIT_36(256'h2000000079000000D2000000C60000004B0000003E00000056000000FC000000),
   .INIT_37(256'hF40000005A000000CD00000078000000FE000000C0000000DB0000009A000000),
   .INIT_38(256'h31000000C7000000070000008800000033000000A8000000DD0000001F000000),
   .INIT_39(256'h5F000000EC0000008000000027000000590000001000000012000000B1000000),
   .INIT_3A(256'h0D0000004A000000B500000019000000A90000007F0000005100000060000000),
   .INIT_3B(256'hEF0000009C000000C9000000930000009F0000007A000000E50000002D000000),
   .INIT_3C(256'hB0000000F50000002A000000AE0000004D0000003B000000E0000000A0000000),
   .INIT_3D(256'h610000009900000053000000830000003C000000BB000000EB000000C8000000),
   .INIT_3E(256'h26000000D600000077000000BA0000007E000000040000002B00000017000000),
   .INIT_3F(256'h7D0000000C0000002100000055000000630000001400000069000000E1000000),
   // TABLE T2 (t_in)
   .INIT_40(256'h03934BE358ABACFA45F11F9D6BCB3BAB5E963A27A4C31A1765537E41A75051F4),
   .INIT_41(256'hA38FB56244802635CBD7C52AD7FC4FE54C25F502769188CC6DF6AD76FA552030),
   .INIT_42(256'hF9C66BD397A38D46F012814C7502C32FC0E15DFE0E9845EA1B6725BA5A49DEB1),
   .INIT_43(256'hC8448EC9692949E021D35874832DD4BE59DA95527AEBBF6D9C9515925FE7038F),
   .INIT_44(256'h3AB47DCEAC66C920AD17F0884FB6BEE171DD27B93E6B99587978F48E896A75C2),
   .INIT_45(256'h2B94F908A01CFE81AE84BB6B77E0B1647F456253336097513182E51A4A1863DF),
   .INIT_46(256'hAB2A66558F57E31F02E2724BD323AB73F8B7527B6C8794DEFD198F4568587048),
   .INIT_47(256'h825CED166ABA0203A5B223BF87F2302808A5D3377B9A86C5C2032FB52807B2EB),
   .INIT_48(256'hFE8AC4A6621FD134BED50605F4CD65DAE2A14E69F2F0F307B492A7791C2B8ACF),
   .INIT_49(256'h1051BD6E9F065E71EFAA4060EC390B83EB75A4F6E132058A55A0A2F3539D342E),
   .INIT_4A(256'h15FF6050D46F04065D0571C48DB59154BD464DE605AEDD3E063D96DD8AF93E21),
   .INIT_4B(256'hEEDB79C85B38E7198B88078942BDB0E89E7767D943CC8940E997D6BDFB241998),
   .INIT_4C(256'h724E6C5A70AC1E11ED48322B86830980000000001EC9F8840FE97C420A47A17C),
   .INIT_4D(256'h2E3A243654D19B5BA621685CD9640A0F3927362DD51E3DAE38560F85FFFBFD0E),
   .INIT_4E(256'h1A161C124B695A7720A261DCC54F80C0919E1B9B96D2B4EEE70F935767B10C0A),
   .INIT_4F(256'hA9C8141EA8B92DB6C7ADF28B0D0B0E09171D121BE0433C222AE5C0A0BA0AE293),
   .INIT_50(256'h7E345BFB3BC54466F5BC5C72269FF70160FDA37FDDBBEE99074CAF75198557F1),
   .INIT_51(256'h112084C62240139785104263DCCAD731F163B8E4FC68B6EDC6DCCB2329768B43),
   .INIT_52(256'hE3D077C152EC0D8630F3DCB22F4B1D9EA16DC7293211AEF93DF8D2BB247D854A),
   .INIT_53(256'h90EF22332CD8567D3F1AA0F08CC4A8FC642247E948FA1194B999A970166C2BB3),
   .INIT_54(256'hBFA43FAD8E26DAB7DE28A57A81CFA6F50B3698D4A2FE8CCAD1C1D9384EC78749),
   .INIT_55(256'hAFF582C3F75E2E39B8E890D813C2F68D4662547ECC9B6A5F920D50789DE42C3A),
   .INIT_56(256'hBB7BDB3B636EE89C7DA71018993BC8AC12B3CF252DA96FD5937C69D080BE9F5D),
   .INIT_57(256'hE8E6EF15CF0821BCE67EAAFF6E65E6959AA8834FB701EC9A18F46E597809CD26),
   .INIT_58(256'h66C035A29430C6A523312A3FB2AF31A47CD629B009D4EA9F36CE4A6F9BD9BAE7),
   .INIT_59(256'hF62F1791500E7FCDDAF741EC984AF104D81533A7D0B0E090CAA6FC82BC37744E),
   .INIT_5A(256'h517F46651FB8C12C881B4C6AB5E39ED104DFE4964D54CCAAB04D43EFD68D764D),
   .INIT_5B(256'h47136DD65633E910D25292DB1D5AB367412EFB0B7473FA87355D018CEA049D5E),
   .INIT_5C(256'hB13C7A47E5EDE11CC935B76127EECEA93C89EB13148E59F80C7A37A1618C9AD7),
   .INIT_5D(256'hDB8678446F14DF3DAA5B5FFDCDEA53F737BF73C7CE791814733F55F2DF599CD2),
   .INIT_5E(256'h9541FF0D498B283C250CBCE2C372161D405FC2A3342C3824C43EB968F381CAAF),
   .INIT_5F(256'h5742D0B85C74486CB670D53284617BCBC1906456E49CD8B4B3DE080C017139A8),
   // TABLE T2 (t_il)
   .INIT_60(256'h000038000000A50000003600000030000000D50000006A000000090000005200),
   .INIT_61(256'h0000FB000000D7000000F3000000810000009E000000A300000040000000BF00),
   .INIT_62(256'h000087000000FF0000002F0000009B0000008200000039000000E30000007C00),
   .INIT_63(256'h0000CB000000E9000000DE000000C400000044000000430000008E0000003400),
   .INIT_64(256'h00003D00000023000000C2000000A600000032000000940000007B0000005400),
   .INIT_65(256'h00004E000000C3000000FA000000420000000B000000950000004C000000EE00),
   .INIT_66(256'h0000B200000024000000D90000002800000066000000A10000002E0000000800),
   .INIT_67(256'h000025000000D10000008B0000006D00000049000000A20000005B0000007600),
   .INIT_68(256'h00001600000098000000680000008600000064000000F6000000F80000007200),
   .INIT_69(256'h000092000000B6000000650000005D000000CC0000005C000000A4000000D400),
   .INIT_6A(256'h0000DA000000B9000000ED000000FD0000005000000048000000700000006C00),
   .INIT_6B(256'h0000840000009D0000008D000000A70000005700000046000000150000005E00),
   .INIT_6C(256'h00000A000000D3000000BC0000008C00000000000000AB000000D80000009000),
   .INIT_6D(256'h00000600000045000000B3000000B80000000500000058000000E4000000F700),
   .INIT_6E(256'h0000020000000F0000003F000000CA0000008F0000001E0000002C000000D000),
   .INIT_6F(256'h00006B0000008A000000130000000100000003000000BD000000AF000000C100),
   .INIT_70(256'h0000EA000000DC000000670000004F0000004100000011000000910000003A00),
   .INIT_71(256'h000073000000E6000000B4000000F0000000CE000000CF000000F20000009700),
   .INIT_72(256'h00008500000035000000AD000000E70000002200000074000000AC0000009600),
   .INIT_73(256'h00006E000000DF000000750000001C000000E800000037000000F9000000E200),
   .INIT_74(256'h000089000000C5000000290000001D000000710000001A000000F10000004700),
   .INIT_75(256'h00001B000000BE00000018000000AA0000000E00000062000000B70000006F00),
   .INIT_76(256'h00002000000079000000D2000000C60000004B0000003E00000056000000FC00),
   .INIT_77(256'h0000F40000005A000000CD00000078000000FE000000C0000000DB0000009A00),
   .INIT_78(256'h000031000000C7000000070000008800000033000000A8000000DD0000001F00),
   .INIT_79(256'h00005F000000EC0000008000000027000000590000001000000012000000B100),
   .INIT_7A(256'h00000D0000004A000000B500000019000000A90000007F000000510000006000),
   .INIT_7B(256'h0000EF0000009C000000C9000000930000009F0000007A000000E50000002D00),
   .INIT_7C(256'h0000B0000000F50000002A000000AE0000004D0000003B000000E0000000A000),
   .INIT_7D(256'h0000610000009900000053000000830000003C000000BB000000EB000000C800),
   .INIT_7E(256'h000026000000D600000077000000BA0000007E000000040000002B0000001700),
   .INIT_7F(256'h00007D0000000C0000002100000055000000630000001400000069000000E100),	
    // The next set of INITP_xx are f6743000000000000000or the parity bits
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)) 
	
	RAMB36_0 (
    .CASCADEOUTLATA(             ), // 1-bit cascade A latch output
    .CASCADEOUTLATB(             ), // 1-bit cascade B latch output
    .CASCADEOUTREGA(             ), // 1-bit cascade A register output
    .CASCADEOUTREGB(             ), // 1-bit cascade B register output
    .DOA           (bram0a_data  ), // 32-bit A port data output
    .DOB           (bram0b_data  ), // 32-bit B port data output
    .DOPA          (             ), // 4-bit A port parity data output
    .DOPB          (             ), // 4-bit B port parity data output
    .ADDRA         (bram0a_addr  ), // 16-bit A port address input
    .ADDRB         (bram0b_addr  ), // 16-bit B port address input
    .CASCADEINLATA (1'b0         ), // 1-bit cascade A latch input
    .CASCADEINLATB (1'b0         ), // 1-bit cascade B latch input
    .CASCADEINREGA (1'b0         ), // 1-bit cascade A register input
    .CASCADEINREGB (1'b0         ), // 1-bit cascade B register input
    .CLKA          (CLK          ), // 1-bit A port clock input
    .CLKB          (CLK          ), // 1-bit B port clock input
    .DIA           (32'd0        ), // 32-bit A port data input
    .DIB           (32'd0        ), // 32-bit B port data input
    .DIPA          (4'd0         ), // 4-bit A port parity data input
    .DIPB          (4'd0         ), // 4-bit B port parity data input
    .ENA           (1'b1         ), // 1-bit A port enable input
    .ENB           (1'b1         ), // 1-bit B port enable input
    .REGCEA        (1'b1         ), // 1-bit A port register enable input
    .REGCEB        (1'b1         ), // 1-bit B port register enable input
    .SSRA          (1'b0         ), // 1-bit A port set/reset input
    .SSRB          (1'b0         ), // 1-bit B port set/reset input
    .WEA           (4'd0         ), // 4-bit A port write enable input
    .WEB           (4'd0         )  // 4-bit B port write enable input
  );

    // shift control for column 0 and 1  
  always @(posedge CLK) begin
    if (TSH[3]) bram0a_data_p <= {bram0a_data[07:00], bram0a_data[31:08]};
    else        bram0a_data_p <= bram0a_data;
    if (TSH[2]) bram0b_data_p <= {bram0b_data[07:00], bram0b_data[31:08]};
    else        bram0b_data_p <= bram0b_data;
  end

  // control input to A:B input of column 0's DSP
  assign dsp0a_din = POB ? PTX : bram0a_data_p;
  
  DSP48E #(
    .ACASCREG                       (1               ), // Number of pipeline registers between A/ACIN input and ACOUT output, 0, 1, or 2
    .ALUMODEREG                     (0               ), // Number of pipeline registers on ALUMODE input, 0 or 1
    .AREG                           (1               ), // Number of pipeline registers on the A input, 0, 1 or 2
    .AUTORESET_PATTERN_DETECT       ("FALSE"         ), // Auto-reset upon pattern detect, "TRUE" or "FALSE"
    .AUTORESET_PATTERN_DETECT_OPTINV("MATCH"         ), // Reset if "MATCH" or "NOMATCH"
    .A_INPUT                        ("DIRECT"        ), // Selects A input used, "DIRECT" (A port) or "CASCADE" (ACIN port)
    .BCASCREG                       (1               ), // Number of pipeline registers between B/BCIN input and BCOUT output, 0, 1, or 2
    .BREG                           (1               ), // Number of pipeline registers on the B input, 0, 1 or 2
    .B_INPUT                        ("DIRECT"        ), // Selects B input used, "DIRECT" (B port) or "CASCADE" (BCIN port)
    .CARRYINREG                     (0               ), // Number of pipeline registers for the CARRYIN input, 0 or 1
    .CARRYINSELREG                  (0               ), // Number of pipeline registers for the CARRYINSEL input, 0 or 1
    .CREG                           (1               ), // Number of pipeline registers on the C input, 0 or 1
    .MASK                           (48'h3fffffffffff), // 48-bit Mask value for pattern detect
    .MREG                           (0               ), // Number of multiplier pipeline registers, 0 or 1
    .MULTCARRYINREG                 (0               ), // Number of pipeline registers for multiplier carry in bit, 0 or 1
    .OPMODEREG                      (1               ), // Number of pipeline registers on OPMODE input, 0 or 1
    .PATTERN                        (48'h000000000000), // 48-bit Pattern match for pattern detect
    .PREG                           (1               ), // Number of pipeline registers on the P output, 0 or 1
    .SEL_MASK                       ("MASK"          ), // Select mask value between the "MASK" value or the value on the "C" port
    .SEL_PATTERN                    ("PATTERN"       ), // Select pattern value between the "PATTERN" value or the value on the "C" port
    .SEL_ROUNDING_MASK              ("SEL_MASK"      ), // "SEL_MASK", "MODE1", "MODE2"
    .USE_MULT                       ("NONE"          ), // Select multiplier usage, "MULT" (MREG => 0), "MULT_S" (MREG => 1), "NONE" (no multiplier)
    .USE_PATTERN_DETECT             ("NO_PATDET"     ), // Enable pattern detect, "PATDET", "NO_PATDET"
    .USE_SIMD                       ("ONE48"         ))  // SIMD selection, "ONE48", "TWO24", "FOUR12"
  DSP48E_0a (
    .ACOUT         (                  ), // 30-bit A port cascade output
    .BCOUT         (                  ), // 18-bit B port cascade output
    .CARRYCASCOUT  (                  ), // 1-bit cascade carry output
    .CARRYOUT      (                  ), // 4-bit carry output
    .MULTSIGNOUT   (                  ), // 1-bit multiplier sign cascade output
    .OVERFLOW      (                  ), // 1-bit overflow in add/acc output
    .P             (                  ), // 48-bit output
    .PATTERNBDETECT(                  ), // 1-bit active high pattern bar detect output
    .PATTERNDETECT (                  ), // 1-bit active high pattern detect output
    .PCOUT         (dsp0a_pdata       ), // 48-bit cascade output
    .UNDERFLOW     (                  ), // 1-bit active high underflow in add/acc output
    .A             ({16'd0,dsp0a_din[31:18]}), // 30-bit A data input
    .ACIN          (                  ), // 30-bit A cascade data input
    .ALUMODE       (4'b0100           ), // 4-bit ALU control input
    .B             (dsp0a_din[17:00]  ), // 18-bit B data input
    .BCIN          (                  ), // 18-bit B cascade input
    .C             ({16'd0,KEY}       ), // 48-bit C data input
    .CARRYCASCIN   (                  ), // 1-bit cascade carry input
    .CARRYIN       (                  ), // 1-bit carry input signal
    .CARRYINSEL    (                  ), // 3-bit carry select input
    .CEA1          (1'b0              ), // 1-bit active high clock enable input for 1st stage A registers
    .CEA2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage A registers
    .CEALUMODE     (1'b0              ), // 1-bit active high clock enable input for ALUMODE registers
    .CEB1          (1'b0              ), // 1-bit active high clock enable input for 1st stage B registers
    .CEB2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage B registers
    .CEC           (1'b1              ), // 1-bit active high clock enable input for C registers
    .CECARRYIN     (1'b0              ), // 1-bit active high clock enable input for CARRYIN register
    .CECTRL        (1'b1              ), // 1-bit active high clock enable input for OPMODE and carry registers
    .CEM           (1'b0              ), // 1-bit active high clock enable input for multiplier registers
    .CEMULTCARRYIN (1'b0              ), // 1-bit active high clock enable for multiplier carry in register
    .CEP           (1'b1              ), // 1-bit active high clock enable input for P registers
    .CLK           (CLK               ), // Clock input
    .MULTSIGNIN    (                  ), // 1-bit multiplier sign input
    .OPMODE        (C_XOR_AB          ), // 7-bit operation mode input
    .PCIN          (                  ), // 48-bit P cascade input
    .RSTA          (1'b0              ), // 1-bit reset input for A pipeline registers
    .RSTALLCARRYIN (1'b0              ), // 1-bit reset input for carry pipeline registers
    .RSTALUMODE    (1'b0              ), // 1-bit reset input for ALUMODE pipeline registers
    .RSTB          (1'b0              ), // 1-bit reset input for B pipeline registers
    .RSTC          (1'b0              ), // 1-bit reset input for C pipeline registers
    .RSTCTRL       (1'b0              ), // 1-bit reset input for OPMODE pipeline registers
    .RSTM          (1'b0              ), // 1-bit reset input for multiplier registers
    .RSTP          (1'b0              ) // 1-bit reset input for P pipeline registers
  );

  DSP48E #(
    .ACASCREG                       (1               ), // Number of pipeline registers between A/ACIN input and ACOUT output, 0, 1, or 2
    .ALUMODEREG                     (0               ), // Number of pipeline registers on ALUMODE input, 0 or 1
    .AREG                           (1               ), // Number of pipeline registers on the A input, 0, 1 or 2
    .AUTORESET_PATTERN_DETECT       ("FALSE"         ), // Auto-reset upon pattern detect, "TRUE" or "FALSE"
    .AUTORESET_PATTERN_DETECT_OPTINV("MATCH"         ), // Reset if "MATCH" or "NOMATCH"
    .A_INPUT                        ("DIRECT"        ), // Selects A input used, "DIRECT" (A port) or "CASCADE" (ACIN port)
    .BCASCREG                       (1               ), // Number of pipeline registers between B/BCIN input and BCOUT output, 0, 1, or 2
    .BREG                           (1               ), // Number of pipeline registers on the B input, 0, 1 or 2
    .B_INPUT                        ("DIRECT"        ), // Selects B input used, "DIRECT" (B port) or "CASCADE" (BCIN port)
    .CARRYINREG                     (0               ), // Number of pipeline registers for the CARRYIN input, 0 or 1
    .CARRYINSELREG                  (0               ), // Number of pipeline registers for the CARRYINSEL input, 0 or 1
    .CREG                           (1               ), // Number of pipeline registers on the C input, 0 or 1
    .MASK                           (48'h3fffffffffff), // 48-bit Mask value for pattern detect
    .MREG                           (0               ), // Number of multiplier pipeline registers, 0 or 1
    .MULTCARRYINREG                 (0               ), // Number of pipeline registers for multiplier carry in bit, 0 or 1
    .OPMODEREG                      (1               ), // Number of pipeline registers on OPMODE input, 0 or 1
    .PATTERN                        (48'h000000000000), // 48-bit Pattern match for pattern detect
    .PREG                           (1               ), // Number of pipeline registers on the P output, 0 or 1
    .SEL_MASK                       ("MASK"          ), // Select mask value between the "MASK" value or the value on the "C" port
    .SEL_PATTERN                    ("PATTERN"       ), // Select pattern value between the "PATTERN" value or the value on the "C" port
    .SEL_ROUNDING_MASK              ("SEL_MASK"      ), // "SEL_MASK", "MODE1", "MODE2"
    .USE_MULT                       ("NONE"          ), // Select multiplier usage, "MULT" (MREG => 0), "MULT_S" (MREG => 1), "NONE" (no multiplier)
    .USE_PATTERN_DETECT             ("NO_PATDET"     ), // Enable pattern detect, "PATDET", "NO_PATDET"
    .USE_SIMD                       ("ONE48"         )) // SIMD selection, "ONE48", "TWO24", "FOUR12"
  DSP48E_0b (
    .ACOUT         (                  ), // 30-bit A port cascade output
    .BCOUT         (                  ), // 18-bit B port cascade output
    .CARRYCASCOUT  (                  ), // 1-bit cascade carry output
    .CARRYOUT      (                  ), // 4-bit carry output
    .MULTSIGNOUT   (                  ), // 1-bit multiplier sign cascade output
    .OVERFLOW      (                  ), // 1-bit overflow in add/acc output
    .P             (                  ), // 48-bit output
    .PATTERNBDETECT(                  ), // 1-bit active high pattern bar detect output
    .PATTERNDETECT (                  ), // 1-bit active high pattern detect output
    .PCOUT         (dsp0b_pdata       ), // 48-bit cascade output
    .UNDERFLOW     (                  ), // 1-bit active high underflow in add/acc output
    .A             ({16'd0,bram0b_data_p[31:18]}), // 30-bit A data input
    .ACIN          (                  ), // 30-bit A cascade data input
    .ALUMODE       (4'b0100           ), // 4-bit ALU control input
    .B             (bram0b_data_p[17:00]), // 18-bit B data input
    .BCIN          (                  ), // 18-bit B cascade input
    .C             ({16'd0,KEY}       ), // 48-bit C data input
    .CARRYCASCIN   (                  ), // 1-bit cascade carry input
    .CARRYIN       (                  ), // 1-bit carry input signal
    .CARRYINSEL    (                  ), // 3-bit carry select input
    .CEA1          (1'b0              ), // 1-bit active high clock enable input for 1st stage A registers
    .CEA2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage A registers
    .CEALUMODE     (1'b0              ), // 1-bit active high clock enable input for ALUMODE registers
    .CEB1          (1'b0              ), // 1-bit active high clock enable input for 1st stage B registers
    .CEB2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage B registers
    .CEC           (1'b1              ), // 1-bit active high clock enable input for C registers
    .CECARRYIN     (1'b0              ), // 1-bit active high clock enable input for CARRYIN register
    .CECTRL        (1'b1              ), // 1-bit active high clock enable input for OPMODE and carry registers
    .CEM           (1'b0              ), // 1-bit active high clock enable input for multiplier registers
    .CEMULTCARRYIN (1'b0              ), // 1-bit active high clock enable for multiplier carry in register
    .CEP           (1'b1              ), // 1-bit active high clock enable input for P registers
    .CLK           (CLK               ), // Clock input
    .MULTSIGNIN    (                  ), // 1-bit multiplier sign input
    .OPMODE        (PCIN_XOR_AB       ), // 7-bit operation mode input
    .PCIN          (dsp0a_pdata       ), // 48-bit P cascade input
    .RSTA          (RXR[2]            ), // 1-bit reset input for A pipeline registers
    .RSTALLCARRYIN (1'b0              ), // 1-bit reset input for carry pipeline registers
    .RSTALUMODE    (1'b0              ), // 1-bit reset input for ALUMODE pipeline registers
    .RSTB          (RXR[2]            ), // 1-bit reset input for B pipeline registers
    .RSTC          (1'b0              ), // 1-bit reset input for C pipeline registers
    .RSTCTRL       (1'b0              ), // 1-bit reset input for OPMODE pipeline registers
    .RSTM          (1'b0              ), // 1-bit reset input for multiplier registers
    .RSTP          (1'b0              ) // 1-bit reset input for P pipeline registers
  );

  RAMB36 #(
    .DOA_REG            (1            ), // Optional output registers on A port (0 or 1)
    .DOB_REG            (1            ), // Optional output registers on B port (0 or 1)
    .INIT_A             (36'h000000000), // Initial values on A output port
    .INIT_B             (36'h000000000), // Initial values on B output port
    .RAM_EXTENSION_A    ("NONE"       ), // "UPPER", "LOWER" or "NONE" when cascaded
    .RAM_EXTENSION_B    ("NONE"       ), // "UPPER", "LOWER" or "NONE" when cascaded
    .READ_WIDTH_A       (36           ), // Valid values are 1, 2, 4, 9, 18, or 36
    .READ_WIDTH_B       (36           ), // Valid values are 1, 2, 4, 9, 18, or 36
    .SIM_COLLISION_CHECK("NONE"       ), // Collision check enable "ALL", "WARNING_ONLY", "GENERATE_X_ONLY" or "NONE"
    .SRVAL_A            (36'h000000000), // Set/Reset value for A port output
    .SRVAL_B            (36'h000000000), // Set/Reset value for B port output
    .WRITE_MODE_A       ("READ_FIRST" ), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
    .WRITE_MODE_B       ("READ_FIRST" ), // "WRITE_FIRST", "READ_FIRST", or "NO_CHANGE"
    .WRITE_WIDTH_A      (36           ), // Valid values are 1, 2, 4, 9, 18, or 36
    .WRITE_WIDTH_B      (36           ), // Valid values are 1, 2, 4, 9, 18, or 36

   // TABLE T0 (t_in)
   .INIT_00(256'h4BE30393ACFA58AB1F9D45F13BAB6BCB3A275E961A17A4C37E41655351F4A750),
   .INIT_01(256'hB562A38F26354480C52ACBD74FE5D7FCF5024C2588CC7691AD766DF62030FA55),
   .INIT_02(256'h6BD3F9C68D4697A3814CF012C32F75025DFEC0E145EA0E9825BA1B67DEB15A49),
   .INIT_03(256'h8EC9C84449E06929587421D3D4BE832D955259DABF6D7AEB15929C95038F5FE7),
   .INIT_04(256'h7DCE3AB4C920AC66F088AD17BEE14FB627B971DD99583E6BF48E797875C2896A),
   .INIT_05(256'hF9082B94FE81A01CBB6BAE84B16477E062537F4597513360E51A318263DF4A18),
   .INIT_06(256'h6655AB2AE31F8F57724B02E2AB73D323527BF8B794DE6C878F45FD1970486858),
   .INIT_07(256'hED16825C02036ABA23BFA5B2302887F2D33708A586C57B9A2FB5C203B2EB2807),
   .INIT_08(256'hC4A6FE8AD134621F0605BED565DAF4CD4E69E2A1F307F2F0A779B4928ACF1C2B),
   .INIT_09(256'hBD6E10515E719F064060EFAA0B83EC39A4F6EB75058AE132A2F355A0342E539D),
   .INIT_0A(256'h605015FF0406D46F71C45D0591548DB54DE6BD46DD3E05AE96DD063D3E218AF9),
   .INIT_0B(256'h79C8EEDBE7195B3807898B88B0E842BD67D99E77894043CCD6BDE9971998FB24),
   .INIT_0C(256'h6C5A724E1E1170AC322BED480980868300000000F8841EC97C420FE9A17C0A47),
   .INIT_0D(256'h24362E3A9B5B54D1685CA6210A0FD964362D39273DAED51E0F853856FD0EFFFB),
   .INIT_0E(256'h1C121A165A774B6961DC20A280C0C54F1B9B919EB4EE96D29357E70F0C0A67B1),
   .INIT_0F(256'h141EA9C82DB6A8B9F28BC7AD0E090D0B121B171D3C22E043C0A02AE5E293BA0A),
   .INIT_10(256'h5BFB7E3444663BC55C72F5BCF701269FA37F60FDEE99DDBBAF75074C57F11985),
   .INIT_11(256'h84C611201397224042638510D731DCCAB8E4F163B6EDFC68CB23C6DC8B432976),
   .INIT_12(256'h77C1E3D00D8652ECDCB230F31D9E2F4BC729A16DAEF93211D2BB3DF8854A247D),
   .INIT_13(256'h223390EF567D2CD8A0F03F1AA8FC8CC447E96422119448FAA970B9992BB3166C),
   .INIT_14(256'h3FADBFA4DAB78E26A57ADE28A6F581CF98D40B368CCAA2FED938D1C187494EC7),
   .INIT_15(256'h82C3AFF52E39F75E90D8B8E8F68D13C2547E46626A5FCC9B5078920D2C3A9DE4),
   .INIT_16(256'hDB3BBB7BE89C636E10187DA7C8AC993BCF2512B36FD52DA969D0937C9F5D80BE),
   .INIT_17(256'hEF15E8E621BCCF08AAFFE67EE6956E65834F9AA8EC9AB7016E5918F4CD267809),
   .INIT_18(256'h35A266C0C6A594302A3F233131A4B2AF29B07CD6EA9F09D44A6F36CEBAE79BD9),
   .INIT_19(256'h1791F62F7FCD500E41ECDAF7F104984A33A7D815E090D0B0FC82CAA6744EBC37),
   .INIT_1A(256'h4665517FC12C1FB84C6A881B9ED1B5E3E49604DFCCAA4D5443EFB04D764DD68D),
   .INIT_1B(256'h6DD64713E910563392DBD252B3671D5AFB0B412EFA877473018C355D9D5EEA04),
   .INIT_1C(256'h7A47B13CE11CE5EDB761C935CEA927EEEB133C8959F8148E37A10C7A9AD7618C),
   .INIT_1D(256'h7844DB86DF3D6F145FFDAA5B53F7CDEA73C737BF1814CE7955F2733F9CD2DF59),
   .INIT_1E(256'hFF0D9541283C498BBCE2250C161DC372C2A3405F3824342CB968C43ECAAFF381),
   .INIT_1F(256'hD0B85742486C5C74D532B6707BCB84616456C190D8B4E49C080CB3DE39A80171),
   // TABLE T0 (t_il)
   .INIT_20(256'h38000000A50000003600000030000000D50000006A0000000900000052000000),
   .INIT_21(256'hFB000000D7000000F3000000810000009E000000A300000040000000BF000000),
   .INIT_22(256'h87000000FF0000002F0000009B0000008200000039000000E30000007C000000),
   .INIT_23(256'hCB000000E9000000DE000000C400000044000000430000008E00000034000000),
   .INIT_24(256'h3D00000023000000C2000000A600000032000000940000007B00000054000000),
   .INIT_25(256'h4E000000C3000000FA000000420000000B000000950000004C000000EE000000),
   .INIT_26(256'hB200000024000000D90000002800000066000000A10000002E00000008000000),
   .INIT_27(256'h25000000D10000008B0000006D00000049000000A20000005B00000076000000),
   .INIT_28(256'h1600000098000000680000008600000064000000F6000000F800000072000000),
   .INIT_29(256'h92000000B6000000650000005D000000CC0000005C000000A4000000D4000000),
   .INIT_2A(256'hDA000000B9000000ED000000FD0000005000000048000000700000006C000000),
   .INIT_2B(256'h840000009D0000008D000000A70000005700000046000000150000005E000000),
   .INIT_2C(256'h0A000000D3000000BC0000008C00000000000000AB000000D800000090000000),
   .INIT_2D(256'h0600000045000000B3000000B80000000500000058000000E4000000F7000000),
   .INIT_2E(256'h020000000F0000003F000000CA0000008F0000001E0000002C000000D0000000),
   .INIT_2F(256'h6B0000008A000000130000000100000003000000BD000000AF000000C1000000),
   .INIT_30(256'hEA000000DC000000670000004F0000004100000011000000910000003A000000),
   .INIT_31(256'h73000000E6000000B4000000F0000000CE000000CF000000F200000097000000),
   .INIT_32(256'h8500000035000000AD000000E70000002200000074000000AC00000096000000),
   .INIT_33(256'h6E000000DF000000750000001C000000E800000037000000F9000000E2000000),
   .INIT_34(256'h89000000C5000000290000001D000000710000001A000000F100000047000000),
   .INIT_35(256'h1B000000BE00000018000000AA0000000E00000062000000B70000006F000000),
   .INIT_36(256'h2000000079000000D2000000C60000004B0000003E00000056000000FC000000),
   .INIT_37(256'hF40000005A000000CD00000078000000FE000000C0000000DB0000009A000000),
   .INIT_38(256'h31000000C7000000070000008800000033000000A8000000DD0000001F000000),
   .INIT_39(256'h5F000000EC0000008000000027000000590000001000000012000000B1000000),
   .INIT_3A(256'h0D0000004A000000B500000019000000A90000007F0000005100000060000000),
   .INIT_3B(256'hEF0000009C000000C9000000930000009F0000007A000000E50000002D000000),
   .INIT_3C(256'hB0000000F50000002A000000AE0000004D0000003B000000E0000000A0000000),
   .INIT_3D(256'h610000009900000053000000830000003C000000BB000000EB000000C8000000),
   .INIT_3E(256'h26000000D600000077000000BA0000007E000000040000002B00000017000000),
   .INIT_3F(256'h7D0000000C0000002100000055000000630000001400000069000000E1000000),
   // TABLE T2 (t_in)
   .INIT_40(256'h03934BE358ABACFA45F11F9D6BCB3BAB5E963A27A4C31A1765537E41A75051F4),
   .INIT_41(256'hA38FB56244802635CBD7C52AD7FC4FE54C25F502769188CC6DF6AD76FA552030),
   .INIT_42(256'hF9C66BD397A38D46F012814C7502C32FC0E15DFE0E9845EA1B6725BA5A49DEB1),
   .INIT_43(256'hC8448EC9692949E021D35874832DD4BE59DA95527AEBBF6D9C9515925FE7038F),
   .INIT_44(256'h3AB47DCEAC66C920AD17F0884FB6BEE171DD27B93E6B99587978F48E896A75C2),
   .INIT_45(256'h2B94F908A01CFE81AE84BB6B77E0B1647F456253336097513182E51A4A1863DF),
   .INIT_46(256'hAB2A66558F57E31F02E2724BD323AB73F8B7527B6C8794DEFD198F4568587048),
   .INIT_47(256'h825CED166ABA0203A5B223BF87F2302808A5D3377B9A86C5C2032FB52807B2EB),
   .INIT_48(256'hFE8AC4A6621FD134BED50605F4CD65DAE2A14E69F2F0F307B492A7791C2B8ACF),
   .INIT_49(256'h1051BD6E9F065E71EFAA4060EC390B83EB75A4F6E132058A55A0A2F3539D342E),
   .INIT_4A(256'h15FF6050D46F04065D0571C48DB59154BD464DE605AEDD3E063D96DD8AF93E21),
   .INIT_4B(256'hEEDB79C85B38E7198B88078942BDB0E89E7767D943CC8940E997D6BDFB241998),
   .INIT_4C(256'h724E6C5A70AC1E11ED48322B86830980000000001EC9F8840FE97C420A47A17C),
   .INIT_4D(256'h2E3A243654D19B5BA621685CD9640A0F3927362DD51E3DAE38560F85FFFBFD0E),
   .INIT_4E(256'h1A161C124B695A7720A261DCC54F80C0919E1B9B96D2B4EEE70F935767B10C0A),
   .INIT_4F(256'hA9C8141EA8B92DB6C7ADF28B0D0B0E09171D121BE0433C222AE5C0A0BA0AE293),
   .INIT_50(256'h7E345BFB3BC54466F5BC5C72269FF70160FDA37FDDBBEE99074CAF75198557F1),
   .INIT_51(256'h112084C62240139785104263DCCAD731F163B8E4FC68B6EDC6DCCB2329768B43),
   .INIT_52(256'hE3D077C152EC0D8630F3DCB22F4B1D9EA16DC7293211AEF93DF8D2BB247D854A),
   .INIT_53(256'h90EF22332CD8567D3F1AA0F08CC4A8FC642247E948FA1194B999A970166C2BB3),
   .INIT_54(256'hBFA43FAD8E26DAB7DE28A57A81CFA6F50B3698D4A2FE8CCAD1C1D9384EC78749),
   .INIT_55(256'hAFF582C3F75E2E39B8E890D813C2F68D4662547ECC9B6A5F920D50789DE42C3A),
   .INIT_56(256'hBB7BDB3B636EE89C7DA71018993BC8AC12B3CF252DA96FD5937C69D080BE9F5D),
   .INIT_57(256'hE8E6EF15CF0821BCE67EAAFF6E65E6959AA8834FB701EC9A18F46E597809CD26),
   .INIT_58(256'h66C035A29430C6A523312A3FB2AF31A47CD629B009D4EA9F36CE4A6F9BD9BAE7),
   .INIT_59(256'hF62F1791500E7FCDDAF741EC984AF104D81533A7D0B0E090CAA6FC82BC37744E),
   .INIT_5A(256'h517F46651FB8C12C881B4C6AB5E39ED104DFE4964D54CCAAB04D43EFD68D764D),
   .INIT_5B(256'h47136DD65633E910D25292DB1D5AB367412EFB0B7473FA87355D018CEA049D5E),
   .INIT_5C(256'hB13C7A47E5EDE11CC935B76127EECEA93C89EB13148E59F80C7A37A1618C9AD7),
   .INIT_5D(256'hDB8678446F14DF3DAA5B5FFDCDEA53F737BF73C7CE791814733F55F2DF599CD2),
   .INIT_5E(256'h9541FF0D498B283C250CBCE2C372161D405FC2A3342C3824C43EB968F381CAAF),
   .INIT_5F(256'h5742D0B85C74486CB670D53284617BCBC1906456E49CD8B4B3DE080C017139A8),
   // TABLE T2 (t_il)
   .INIT_60(256'h000038000000A50000003600000030000000D50000006A000000090000005200),
   .INIT_61(256'h0000FB000000D7000000F3000000810000009E000000A300000040000000BF00),
   .INIT_62(256'h000087000000FF0000002F0000009B0000008200000039000000E30000007C00),
   .INIT_63(256'h0000CB000000E9000000DE000000C400000044000000430000008E0000003400),
   .INIT_64(256'h00003D00000023000000C2000000A600000032000000940000007B0000005400),
   .INIT_65(256'h00004E000000C3000000FA000000420000000B000000950000004C000000EE00),
   .INIT_66(256'h0000B200000024000000D90000002800000066000000A10000002E0000000800),
   .INIT_67(256'h000025000000D10000008B0000006D00000049000000A20000005B0000007600),
   .INIT_68(256'h00001600000098000000680000008600000064000000F6000000F80000007200),
   .INIT_69(256'h000092000000B6000000650000005D000000CC0000005C000000A4000000D400),
   .INIT_6A(256'h0000DA000000B9000000ED000000FD0000005000000048000000700000006C00),
   .INIT_6B(256'h0000840000009D0000008D000000A70000005700000046000000150000005E00),
   .INIT_6C(256'h00000A000000D3000000BC0000008C00000000000000AB000000D80000009000),
   .INIT_6D(256'h00000600000045000000B3000000B80000000500000058000000E4000000F700),
   .INIT_6E(256'h0000020000000F0000003F000000CA0000008F0000001E0000002C000000D000),
   .INIT_6F(256'h00006B0000008A000000130000000100000003000000BD000000AF000000C100),
   .INIT_70(256'h0000EA000000DC000000670000004F0000004100000011000000910000003A00),
   .INIT_71(256'h000073000000E6000000B4000000F0000000CE000000CF000000F20000009700),
   .INIT_72(256'h00008500000035000000AD000000E70000002200000074000000AC0000009600),
   .INIT_73(256'h00006E000000DF000000750000001C000000E800000037000000F9000000E200),
   .INIT_74(256'h000089000000C5000000290000001D000000710000001A000000F10000004700),
   .INIT_75(256'h00001B000000BE00000018000000AA0000000E00000062000000B70000006F00),
   .INIT_76(256'h00002000000079000000D2000000C60000004B0000003E00000056000000FC00),
   .INIT_77(256'h0000F40000005A000000CD00000078000000FE000000C0000000DB0000009A00),
   .INIT_78(256'h000031000000C7000000070000008800000033000000A8000000DD0000001F00),
   .INIT_79(256'h00005F000000EC0000008000000027000000590000001000000012000000B100),
   .INIT_7A(256'h00000D0000004A000000B500000019000000A90000007F000000510000006000),
   .INIT_7B(256'h0000EF0000009C000000C9000000930000009F0000007A000000E50000002D00),
   .INIT_7C(256'h0000B0000000F50000002A000000AE0000004D0000003B000000E0000000A000),
   .INIT_7D(256'h0000610000009900000053000000830000003C000000BB000000EB000000C800),
   .INIT_7E(256'h000026000000D600000077000000BA0000007E000000040000002B0000001700),
   .INIT_7F(256'h00007D0000000C0000002100000055000000630000001400000069000000E100),
    // The next set of INITP_xx are for the parity bits
    .INITP_00(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_01(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_02(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_03(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_04(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_05(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_06(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_07(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_08(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_09(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0A(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0B(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0C(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0D(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0E(256'h0000000000000000000000000000000000000000000000000000000000000000),
    .INITP_0F(256'h0000000000000000000000000000000000000000000000000000000000000000)) 
  RAMB36_1 (
    .CASCADEOUTLATA(             ), // 1-bit cascade A latch output
    .CASCADEOUTLATB(             ), // 1-bit cascade B latch output
    .CASCADEOUTREGA(             ), // 1-bit cascade A register output
    .CASCADEOUTREGB(             ), // 1-bit cascade B register output
    .DOA           (bram1a_data  ), // 32-bit A port data output
    .DOB           (bram1b_data  ), // 32-bit B port data output
    .DOPA          (             ), // 4-bit A port parity data output
    .DOPB          (             ), // 4-bit B port parity data output
    .ADDRA         (bram1a_addr  ), // 16-bit A port address input
    .ADDRB         (bram1b_addr  ), // 16-bit B port address input
    .CASCADEINLATA (             ), // 1-bit cascade A latch input
    .CASCADEINLATB (             ), // 1-bit cascade B latch input
    .CASCADEINREGA (             ), // 1-bit cascade A register input
    .CASCADEINREGB (             ), // 1-bit cascade B register input
    .CLKA          (CLK          ), // 1-bit A port clock input
    .CLKB          (CLK          ), // 1-bit B port clock input
    .DIA           (             ), // 32-bit A port data input
    .DIB           (             ), // 32-bit B port data input
    .DIPA          (             ), // 4-bit A port parity data input
    .DIPB          (             ), // 4-bit B port parity data input
    .ENA           (~RST         ), // 1-bit A port enable input
    .ENB           (~RST         ), // 1-bit B port enable input
    .REGCEA        (1'b1         ), // 1-bit A port register enable input
    .REGCEB        (1'b1         ), // 1-bit B port register enable input
    .SSRA          (1'b0         ), // 1-bit A port set/reset input
    .SSRB          (1'b0         ), // 1-bit B port set/reset input
    .WEA           (4'd0         ), // 4-bit A port write enable input
    .WEB           (4'd0         )  // 4-bit B port write enable input
  );

  // shift control for column 2 and 3  
  always @(posedge CLK) begin
    if (TSH[1]) bram1a_data_p <= {bram1a_data[07:00], bram1a_data[31:08]};
    else        bram1a_data_p <= bram1a_data;
    if (TSH[0]) bram1b_data_p <= {bram1b_data[07:00], bram1b_data[31:08]};
    else        bram1b_data_p <= bram1b_data;
  end
  
  DSP48E #(
    .ACASCREG                       (1                 ), // Number of pipeline registers between A/ACIN input and ACOUT output, 0, 1, or 2
    .ALUMODEREG                     (0                 ), // Number of pipeline registers on ALUMODE input, 0 or 1
    .AREG                           (1                 ), // Number of pipeline registers on the A input, 0, 1 or 2
    .AUTORESET_PATTERN_DETECT       ("FALSE"           ), // Auto-reset upon pattern detect, "TRUE" or "FALSE"
    .AUTORESET_PATTERN_DETECT_OPTINV("MATCH"           ), // Reset if "MATCH" or "NOMATCH"
    .A_INPUT                        ("DIRECT"          ), // Selects A input used, "DIRECT" (A port) or "CASCADE" (ACIN port)
    .BCASCREG                       (1                 ), // Number of pipeline registers between B/BCIN input and BCOUT output, 0, 1, or 2
    .BREG                           (1                 ), // Number of pipeline registers on the B input, 0, 1 or 2
    .B_INPUT                        ("DIRECT"          ), // Selects B input used, "DIRECT" (B port) or "CASCADE" (BCIN port)
    .CARRYINREG                     (0                 ), // Number of pipeline registers for the CARRYIN input, 0 or 1
    .CARRYINSELREG                  (0                 ), // Number of pipeline registers for the CARRYINSEL input, 0 or 1
    .CREG                           (1                 ), // Number of pipeline registers on the C input, 0 or 1
    .MASK                           (48'h3fffffffffff  ), // 48-bit Mask value for pattern detect
    .MREG                           (0                 ), // Number of multiplier pipeline registers, 0 or 1
    .MULTCARRYINREG                 (0                 ), // Number of pipeline registers for multiplier carry in bit, 0 or 1
    .OPMODEREG                      (1                 ), // Number of pipeline registers on OPMODE input, 0 or 1
    .PATTERN                        (48'h000000000000  ), // 48-bit Pattern match for pattern detect
    .PREG                           (1                 ), // Number of pipeline registers on the P output, 0 or 1
    .SEL_MASK                       ("MASK"            ), // Select mask value between the "MASK" value or the value on the "C" port
    .SEL_PATTERN                    ("PATTERN"         ), // Select pattern value between the "PATTERN" value or the value on the "C" port
    .SEL_ROUNDING_MASK              ("SEL_MASK"        ), // "SEL_MASK", "MODE1", "MODE2"
    .USE_MULT                       ("NONE"            ), // Select multiplier usage, "MULT" (MREG => 0), "MULT_S" (MREG => 1), "NONE" (no multiplier)
    .USE_PATTERN_DETECT             ("NO_PATDET"       ), // Enable pattern detect, "PATDET", "NO_PATDET"
    .USE_SIMD                       ("ONE48"           )) // SIMD selection, "ONE48", "TWO24", "FOUR12"
  DSP48E_1a (
    .ACOUT         (                  ), // 30-bit A port cascade output
    .BCOUT         (                  ), // 18-bit B port cascade output
    .CARRYCASCOUT  (                  ), // 1-bit cascade carry output
    .CARRYOUT      (                  ), // 4-bit carry output
    .MULTSIGNOUT   (                  ), // 1-bit multiplier sign cascade output
    .OVERFLOW      (                  ), // 1-bit overflow in add/acc output
    .P             (                  ), // 48-bit output
    .PATTERNBDETECT(                  ), // 1-bit active high pattern bar detect output
    .PATTERNDETECT (                  ), // 1-bit active high pattern detect output
    .PCOUT         (dsp1a_pdata       ), // 48-bit cascade output
    .UNDERFLOW     (                  ), // 1-bit active high underflow in add/acc output
    .A             ({16'd0,bram1a_data_p[31:18]}), // 30-bit A data input
    .ACIN          (                  ), // 30-bit A cascade data input
    .ALUMODE       (4'b0100           ), // 4-bit ALU control input
    .B             (bram1a_data_p[17:00]), // 18-bit B data input
    .BCIN          (                  ), // 18-bit B cascade input
    .C             ({16'd0,KEY}       ), // 48-bit C data input
    .CARRYCASCIN   (                  ), // 1-bit cascade carry input
    .CARRYIN       (                  ), // 1-bit carry input signal
    .CARRYINSEL    (                  ), // 3-bit carry select input
    .CEA1          (1'b0              ), // 1-bit active high clock enable input for 1st stage A registers
    .CEA2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage A registers
    .CEALUMODE     (1'b0              ), // 1-bit active high clock enable input for ALUMODE registers
    .CEB1          (1'b0              ), // 1-bit active high clock enable input for 1st stage B registers
    .CEB2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage B registers
    .CEC           (1'b1              ), // 1-bit active high clock enable input for C registers
    .CECARRYIN     (1'b0              ), // 1-bit active high clock enable input for CARRYIN register
    .CECTRL        (1'b1              ), // 1-bit active high clock enable input for OPMODE and carry registers
    .CEM           (1'b0              ), // 1-bit active high clock enable input for multiplier registers
    .CEMULTCARRYIN (1'b0              ), // 1-bit active high clock enable for multiplier carry in register
    .CEP           (1'b1              ), // 1-bit active high clock enable input for P registers
    .CLK           (CLK               ), // Clock input
    .MULTSIGNIN    (                  ), // 1-bit multiplier sign input
    .OPMODE        (PCIN_XOR_AB       ), // 7-bit operation mode input
    .PCIN          (dsp0b_pdata       ), // 48-bit P cascade input
    .RSTA          (RXR[1]            ), // 1-bit reset input for A pipeline registers
    .RSTALLCARRYIN (1'b0              ), // 1-bit reset input for carry pipeline registers
    .RSTALUMODE    (1'b0              ), // 1-bit reset input for ALUMODE pipeline registers
    .RSTB          (RXR[1]            ), // 1-bit reset input for B pipeline registers
    .RSTC          (1'b0              ), // 1-bit reset input for C pipeline registers
    .RSTCTRL       (1'b0              ), // 1-bit reset input for OPMODE pipeline registers
    .RSTM          (1'b0              ), // 1-bit reset input for multiplier registers
    .RSTP          (1'b0              ) // 1-bit reset input for P pipeline registers
  );

  DSP48E #(
    .ACASCREG                       (1               ), // Number of pipeline registers between A/ACIN input and ACOUT output, 0, 1, or 2
    .ALUMODEREG                     (0               ), // Number of pipeline registers on ALUMODE input, 0 or 1
    .AREG                           (1               ), // Number of pipeline registers on the A input, 0, 1 or 2
    .AUTORESET_PATTERN_DETECT       ("FALSE"         ), // Auto-reset upon pattern detect, "TRUE" or "FALSE"
    .AUTORESET_PATTERN_DETECT_OPTINV("MATCH"         ), // Reset if "MATCH" or "NOMATCH"
    .A_INPUT                        ("DIRECT"        ), // Selects A input used, "DIRECT" (A port) or "CASCADE" (ACIN port)
    .BCASCREG                       (1               ), // Number of pipeline registers between B/BCIN input and BCOUT output, 0, 1, or 2
    .BREG                           (1               ), // Number of pipeline registers on the B input, 0, 1 or 2
    .B_INPUT                        ("DIRECT"        ), // Selects B input used, "DIRECT" (B port) or "CASCADE" (BCIN port)
    .CARRYINREG                     (0               ), // Number of pipeline registers for the CARRYIN input, 0 or 1
    .CARRYINSELREG                  (0               ), // Number of pipeline registers for the CARRYINSEL input, 0 or 1
    .CREG                           (1               ), // Number of pipeline registers on the C input, 0 or 1
    .MASK                           (48'h3fffffffffff), // 48-bit Mask value for pattern detect
    .MREG                           (0               ), // Number of multiplier pipeline registers, 0 or 1
    .MULTCARRYINREG                 (0               ), // Number of pipeline registers for multiplier carry in bit, 0 or 1
    .OPMODEREG                      (1               ), // Number of pipeline registers on OPMODE input, 0 or 1
    .PATTERN                        (48'h000000000000), // 48-bit Pattern match for pattern detect
    .PREG                           (1               ), // Number of pipeline registers on the P output, 0 or 1
    .SEL_MASK                       ("MASK"          ), // Select mask value between the "MASK" value or the value on the "C" port
    .SEL_PATTERN                    ("PATTERN"       ), // Select pattern value between the "PATTERN" value or the value on the "C" port
    .SEL_ROUNDING_MASK              ("SEL_MASK"      ), // "SEL_MASK", "MODE1", "MODE2"
    .USE_MULT                       ("NONE"          ), // Select multiplier usage, "MULT" (MREG => 0), "MULT_S" (MREG => 1), "NONE" (no multiplier)
    .USE_PATTERN_DETECT             ("NO_PATDET"     ), // Enable pattern detect, "PATDET", "NO_PATDET"
    .USE_SIMD                       ("ONE48"         )) // SIMD selection, "ONE48", "TWO24", "FOUR12"
  DSP48E_1b (
    .ACOUT         (                  ), // 30-bit A port cascade output
    .BCOUT         (                  ), // 18-bit B port cascade output
    .CARRYCASCOUT  (                  ), // 1-bit cascade carry output
    .CARRYOUT      (                  ), // 4-bit carry output
    .MULTSIGNOUT   (                  ), // 1-bit multiplier sign cascade output
    .OVERFLOW      (                  ), // 1-bit overflow in add/acc output
    .P             (dsp1b_pdata       ), // 48-bit output
    .PATTERNBDETECT(                  ), // 1-bit active high pattern bar detect output
    .PATTERNDETECT (                  ), // 1-bit active high pattern detect output
    .PCOUT         (                  ), // 48-bit cascade output
    .UNDERFLOW     (                  ), // 1-bit active high underflow in add/acc output
    .A             ({16'd0,bram1b_data_p[31:18]}), // 30-bit A data input
    .ACIN          (                  ), // 30-bit A cascade data input
    .ALUMODE       (4'b0100           ), // 4-bit ALU control input
    .B             (bram1b_data_p[17:00]), // 18-bit B data input
    .BCIN          (                  ), // 18-bit B cascade input
    .C             ({16'd0,KEY}       ), // 48-bit C data input
    .CARRYCASCIN   (                  ), // 1-bit cascade carry input
    .CARRYIN       (                  ), // 1-bit carry input signal
    .CARRYINSEL    (                  ), // 3-bit carry select input
    .CEA1          (1'b0              ), // 1-bit active high clock enable input for 1st stage A registers
    .CEA2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage A registers
    .CEALUMODE     (1'b0              ), // 1-bit active high clock enable input for ALUMODE registers
    .CEB1          (1'b0              ), // 1-bit active high clock enable input for 1st stage B registers
    .CEB2          (1'b1              ), // 1-bit active high clock enable input for 2nd stage B registers
    .CEC           (1'b1              ), // 1-bit active high clock enable input for C registers
    .CECARRYIN     (1'b0              ), // 1-bit active high clock enable input for CARRYIN register
    .CECTRL        (1'b1              ), // 1-bit active high clock enable input for OPMODE and carry registers
    .CEM           (1'b0              ), // 1-bit active high clock enable input for multiplier registers
    .CEMULTCARRYIN (1'b0              ), // 1-bit active high clock enable for multiplier carry in register
    .CEP           (1'b1              ), // 1-bit active high clock enable input for P registers
    .CLK           (CLK               ), // Clock input
    .MULTSIGNIN    (                  ), // 1-bit multiplier sign input
    .OPMODE        (PCIN_XOR_AB       ), // 7-bit operation mode input
    .PCIN          (dsp1a_pdata       ), // 48-bit P cascade input
    .RSTA          (RXR[0]            ), // 1-bit reset input for A pipeline registers
    .RSTALLCARRYIN (1'b0              ), // 1-bit reset input for carry pipeline registers
    .RSTALUMODE    (1'b0              ), // 1-bit reset input for ALUMODE pipeline registers
    .RSTB          (RXR[0]            ), // 1-bit reset input for B pipeline registers
    .RSTC          (1'b0              ), // 1-bit reset input for C pipeline registers
    .RSTCTRL       (1'b0              ), // 1-bit reset input for OPMODE pipeline registers
    .RSTM          (1'b0              ), // 1-bit reset input for multiplier registers
    .RSTP          (1'b0              ) // 1-bit reset input for P pipeline registers
  );

endmodule
            